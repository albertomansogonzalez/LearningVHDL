library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity decoder is
	port(	A : in bit_vector (2 downto 0);
		Y : out bit_vector(7 downto 0));
end entity;

architecture arch of decoder is
begin
    with A select
        Y <= "00000001" when "000",
             "00000010" when "001",
             "00000100" when "010",
             "00001000" when "011",
             "00010000" when "100",
             "00100000" when "101",
             "01000000" when "110",
             "10000000" when "111",
             "00000000" when others;
end arch;
